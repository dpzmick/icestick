module spi_slave(
    // fpga signals
    input  clk,
    input  send_in,     // inform that a send be started on `in`. Only valid when `send_avail` is high, must be cleared on next fpga clock
    output send_avail,
    input  [7:0] in,    // when `send_in` is high, in is read and a send is initiated. It is okay to clear `in` on the next `clk`
    output out_avail,   // high when we have something to report reading (the value on `out` will be zero if nothing is being sent)
    output [7:0] out,   // valid value when `out_avail` is high, resets to zero every clock, so get it while its fresh

    // spi signals
    input  SCK,   // Clock generated by the master
    input  SSEL,  // Slave Selection
    input  MOSI,  // Master Out Slave In
    output MISO   // Master In Slave Out
);

// FIXME support reset?

// shift registers to store some spi signals
reg [1:0] sck_  = 2'b0;
reg [1:0] mosi_ = 2'b0;

// temporary storage to push send/recv values into
reg [3:0] send_rem_  = 4'd0;
reg [7:0] sending_   = 8'd0;
reg [3:0] recv_cnt_  = 4'd0;
reg [7:0] receiving_ = 8'd0;

// update shift registers
always @(posedge clk) begin
    if (SSEL) begin
        sck_  <= {sck_[0], SCK};
        mosi_ <= {mosi_[0], MOSI}; // not sure if this needs to be sampled
    end else begin
        sck_      <= 2'b00;
        mosi_     <= 2'b00;
    end
end

// update send and recv buffers
always @(posedge clk) begin
    // if we've finished receiving something recently, "copy" (what's the impact
    // of this) the value, mark it, and reset for next time. This will always
    // run faster than the SPI clock, so it should be fine to "reset" on the
    // fpga clock after the SPI clock that finished producing the value
    // (although that's slow?).

    // Currently letting the counter wrap around, and not clearing anything in
    // `receiving`. By the time we are back to the next `8` in the counter, the
    // entire `receiving` reg will have been cleared anyway.

    if (recv_cnt_ == 4'd8) begin
        out       <= receiving_;
        out_avail <= 1;
    end else begin
        out       <= 8'd0;
        out_avail <= 0;
    end

    if (send_in && send_avail) begin // user wants a send and we have one
        sending_   <= in;
        send_rem_  <= 8;
        send_avail <= 0;
    end else if (send_rem_ == 0) begin // nothing being actively sent
        send_avail <= 1;
    end

    if (SSEL) begin
        if (sck_[1] && !sck_[0]) begin // rising edge, something to sample
            receiving_[7:0] <= {receiving_[6:0], mosi_[1]}; // sampling behind the actual thing will introduce some latency too?
            recv_cnt_       <= recv_cnt_ + 1;

            if (send_rem_ > 0) begin // there's something left for us to send
                MISO      <= sending_[send_rem_-1];
                send_rem_ <= send_rem_ - 1; // should never conflict with the other assignment above? seems bad
            end else begin
                MISO <= 0;
            end
        end
    end
end

endmodule
