module sanity(
    input in,
    output out
);

assign out = ~in;

endmodule
